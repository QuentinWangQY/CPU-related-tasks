library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;  -- ʹ��NUMERIC_STD������з�������

entity ALU is
    port (
        A, B : in STD_LOGIC_VECTOR(31 downto 0);   -- 32λ������
        ALUctr : in STD_LOGIC_VECTOR(2 downto 0);  -- 3λALU�����ź�
        Result : out STD_LOGIC_VECTOR(31 downto 0); -- 32λ������
        Overflow : out STD_LOGIC;                   -- �����־
        Z : out STD_LOGIC                          -- Zero-���־
    );
end ALU;

architecture Behavioral of ALU is
    signal temp_result : STD_LOGIC_VECTOR(31 downto 0);
    signal temp_add, temp_sub : STD_LOGIC_VECTOR(32 downto 0);
    signal overflow_add, overflow_sub : STD_LOGIC;
    signal a_signed, b_signed : SIGNED(31 downto 0);
begin
    -- ����ת��
    a_signed <= SIGNED(A);
    b_signed <= SIGNED(B);
    
    -- �������
    process(A, B, ALUctr, a_signed, b_signed)
    begin
        case ALUctr is
            when "000" => -- ADD: �ӷ�
                temp_result <= A + B;
            when "001" => -- SUB: ����
                temp_result <= A - B;
            when "010" => -- AND: ������
                temp_result <= A and B;
            when "011" => -- OR: ������
                temp_result <= A or B;
            when "100" => -- XOR: �������
                temp_result <= A xor B;
            when "101" => -- NOR: �������
                temp_result <= A nor B;
            when "110" => -- SLT: �з��űȽ� (A < B ? 1 : 0)
                if a_signed < b_signed then
                    temp_result <= X"00000001";
                else
                    temp_result <= X"00000000";
                end if;
            when "111" => -- SLL: �߼����� (B��λλ��)
                temp_result <= STD_LOGIC_VECTOR(SHIFT_LEFT(UNSIGNED(A), to_integer(UNSIGNED(B(4 downto 0)))));
            when others =>
                temp_result <= (others => '0');
        end case;
    end process;
    
    -- ������ (�����з��żӼ���)
    temp_add <= ('0' & A) + ('0' & B);
    temp_sub <= ('0' & A) - ('0' & B);
    
    overflow_add <= '1' when (A(31) = B(31)) and (temp_add(31) /= A(31)) and ALUctr = "000" else '0';
    overflow_sub <= '1' when (A(31) /= B(31)) and (temp_sub(31) /= A(31)) and ALUctr = "001" else '0';
    
    Overflow <= overflow_add or overflow_sub;
    
    -- �����������־
    Result <= temp_result;
    Z <= '1' when temp_result = X"00000000" else '0';
    
end Behavioral;